XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��u��i���b�Mt�ogR��V�mr�����!m�@�@�6 K��N�bj�2,�my�A��#|9t��p�zُ�:m�,&��#a��e'9WI�nj�>*�{�V>G��/�� o�y�7E��N�v\z��E����'�P,S�tݏT�r����7�]�|*�ma\*`!�?�9�S������yb<��Vz���j�Yqm���*���c6L�`G"R�0��0�FP�@�q�W1�8W��ޤ����E�@�SwA��ժb��֕�s?�]��Lb
����C���O)���m��]fb-#(��M��0z1/���/0�L�^HƜ?��c3�\-ؽe�YVZ�5DE�����Ym�lh�|����RmE�I�X�������m���@A��Adw��6�Xz�'e`�'�~���dJ@���}�\�
OB'����������w)")�\D#��K$�@9���}zݴ��H0~'��m�}I��x��V�{e���Y�wP���t�{�PSW��E���'�h�v�S�ԘZoL�#�jD��z7���=��iW��`�M{Pu#�.k�&��G"�C�/�1b�?���`oi|�?<��sp����L�Y���Ȏ�^c�ѹO��a��t�ƋA��~9Hcr�/a�k��+z��nK4o�1�D�Umψm{�B?&�� f��vt�2���nw�[����!�������w�H%�����I�L.R�\	����!����Y��r(�`?<$�S��w��XlxVHYEB    4ba0    1230��-��
�qX���iVg8И��	j�<��#hc��Dxe��?��i*Y�r{>��Ir��Z���N�Ŏ>�/ckR��
��y��z,�i���ٟ.�E�5Zi-x��XSt�Iο��/e�dq�D)1��
�5!��jq�Y$��]I��� }�pt�����-[��?��P.ۆ�`�/g��*�:�)�C�ѷ�D�'��﫬"N�ljǦ1���%������6�����*�r�Дe㤃��мR�1S��e�q�(p�^^MƉ��Z3r9�
Q�g�
l���8I��u���F�%��8�7��y����lk8Š�_��LW�G��� �������C~y�N3�C-r��՝���4-��m�Zʳ"��[d��k�����:9ٴ�,N���@l���:n��;Y6�#Pc=��ݏs�L\�[!�L�������J�q�� I	G��Sf|�Q���^A"�Wp���S���G_ӺL�c^@J���l�v��]W	 K4ᔆ1��]>����D��N]��}�_��a���G ncZ�ϸ�����'�3�(����Yg;�BNAPNY=)g��F�Ś�J9���(�(J�z��f|�K}�k3��|QL����v�������0��p��;C#�����ݽ�/�6�[}�/D�"1����#�fP�B�v�1���H��.����W��@/��sg����/���4ɍ޸/ؾX�F�n��]5�4���p�2Q�`��l���+�H����cn��_��zox50w?o�Ȱ��!�K���!�d�9�<�zg��|gfU��Q�e:D�.�;�����?x%x �b% �Ӏ��lסe+�H��:D<�ķu�p���~Ȼ(�|״0�6�bW���D�2�̖4/*�׬��E�@@����9er6Teּ��`A���l.sx����gʎA-'�;a"}�~|�����\�q�k��i�P��Gd]P�~�zf���|qv5��2q/ʑ�I����#Y/��+ԇU���쐠���"YL(���$��	�s�[T��wf� ��C�x/ˏ���y�P)���9���q�Q-����t'E���냆���=������?g������ͣ����3U���7a�c�KX,/�97i�r�F�/4E�_eF94�����m����5��-2BR��ev�}w�>�?�Cyҡ����sWH��c��}�)�a�[���OM�H����"u�Q�݇�޷E�>�ZY�M�mt��>E���k\��$A �dA��s~�m�SU�i#�9�t��?��[Z��?\�`]�dٓv���V�hs,���fxT�7lg+"�&!o���0��+R�o�B��s��o��5br�Y��q�2�H����{����	�9{>�
�'��XZV�e<�&	�,��-��D�0&r�8LnYhN�N��K%+�N��b��� I��z���������7�}��:�U��{&�3�������V��z���N �s���Ľy�:��0[�`�
�[Ȳ�4$z� E��a�1C�	1y�����6�5�z��8ab�|!2��k=.٬�j~��K��X�a��l�`+�(����8��2�t>�G���'ev
����3���a�NG���q��-����/�{W0����?pE;����j�}*TL�c��C�_@k�C\oA�sK� J�����b^8RXr���J	r�[�����[Qj]����g�b����,����S��6JA!~��F�(���=k��)�}�.������!�A5wng�]hl(�%x��㑲i73��Ur##�/���F�>���0����X<�PHu�k��+E򚙐��N�R?1a�L�ޮj�(y�n���W��!`��L�2������,��
DQ�Oƨ#y�'x�Vc"N�^�J�n��PW��?-d�.����Yf;�O�ѝ�L�^���r]���y��lǲ�:�t���J������b��ڟ~�C�oĻ�R:�w��A�\�X�Q|�K�j*�*A:1��䥋s��'
��l?3�q;��X����A� �\Z�Gd�D�w���Ov�8��+X�O���5�6M��AR��[zo5|<i�G�@�ݲEQ���f���a��^��"@��۵|u��{k� ��mV"qh5��r����Z��倡�qi��n�m�'�o}Q@[c�c�N���q�ˉ�:��Goe4<�jVk��:U��i�Oa%+�Lg7p��:�G��Hh�3��x����]{|��}��=Ŝ��T��F���7��\z���+J�]�X|��O�m	/�d�m�ږU��H?��OPC����;���Qb{�$�Qx�,�,����9��hl�H���Y9o�#��wy�L`�z$��g3�{�N�fZjµɟJi(��c2TkɃ��6���{/�n� ^����tP�"�~H�	����R�r	Y�ᆩ�.s��3�uy�#�?e)V��|�)}r�f�jj��Yd4��tE���{��S],�C	�߹ U]���-���:X���&���Q_)�>$�8 I6�
���}kT *6lg}�wZQ��)���wn�Up�S�yR���r+�i`�kO�����f��g-���Z鰬��Q̕�!#��a3��]�6bw��{rruz�P#���PnIb��U�D �E�"�]�\��g^F2��1�V%�*�D����߮-V;�4.�jҌ��G�<t�`��4�g��L��^���F�_q5�2mZ��9�Cf��Ⱦ=۴I����y���d�L�� �N^�2��%��"����1�l�DZT�Ҳ�]����
g��uD9A�3�)~�������NVBR�b�*�Aڟ���u�wyll�Re�����cLxR
�W��\Q���c�S��r=��߭idw����R�(�ͱ.|�b�6C']��*��x<)��p*g��sG\�aŠ��,�CFc܄�ˉ'&�7����
�B� �@�9�d��/m
�bFk���6֎�iN��ڪ�X���(%�W;��՛U@�1`Q�3�t�l8��%G��r����cH�R�'4�������:I��\8�y�U~��[IK�9�ڝ��i��Q��=�_I$#zl4��f���-=�;�"z�r� (nr���n���w���iA��CɆ���+v�.�n�z�[��m*�^|(�u������\C�� �H��(c�o��]O���{���m��>1�o���J(��,��� � �4K���z��9J� �vЊ&u�r�	()�sl�#���ޮ�ǎr�w�|ʆ�1%��������+��+{ϭ5���BUQ���r��?YK�VW3[�_��,���}sFrv��)�/C���'��	g�0P �+g ��*K㥎�y}V�/K�xE�	��^���B��������������Ԫaoڹ�G��\��������vZ�8�9�t���$�˘}\��}�:Ӽq\6�JUS�����E���o�����pm��/�zW���	����f��`��7�7�}�R�8:����ow)�N,�.6J�}��y���'��\r�G�큢e�{����6TmS�p��e������$�E(����6��
�I}v�]Q�g4�rH��=�W�TZ k�$�ATRˣ�Y���c��ۣ��w_��(��}��e}N=�:��q��ڤ����Ů~�JPjr��g�p�ԛ�m)~.����d^U��u�\qĀt	&�&pZ�u*�����s���k���N��TD�_�@��V��-�I���2��e�)�
;V�������0��͸�"���Ŵ�=�!@a#�/���+}��};Z�MMH��x�윸��}�:ب�k�=$;�"|�	�b�uO����\�fD����[��D�F�rN��{���S�G�K�a)��o��7O闁�BWQ���S�*��b\2�⼑�#�ڃÓuc=<f��t6���M���1�E[�p��~"7����w��#��np�6�U$96�'���A�v�J���ڶf<�؟ݖ?���Wg5������g��&L�d��J	@�VBF6�W^�u��I/Ɗ���9m�أ��N��vN�>~K��z����N��ݫ�z���	�x芒��J}�};%q�Ks��Q S���+T��a����+�iF��&���Fʹ�>�q��� ����;H���+)���S.��l����Q�|�RN��iE`^�EU&�c �YW�(�f��VnZ�uQ��K���a~�7YXv�mƸ�/�HԂ��P�d�`��������7��g�(؉��z>�U�r[�:�.�q/���H���\0ðg���݊O��y�Wb�c���"�޲�Rr�Es�6�������L���Vg?s�����}C���n�u�x[\hQ-\E��P�MZ!+������H����60r7o�Iz������1��#7Mă������
ڎ�7̷dvRI��{z�M����f��>9ZA�Y#%]#�͕iX�f����ݽ�0>�ע�`�x،�8.��T���* ����Nj��J�7�D���~%�X>��Mulu#i�pe����